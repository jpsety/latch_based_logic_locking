// TODO this module should test design
// modes: w/ + w/out scan, locked in parallel, syn, lay
// make a golden model
